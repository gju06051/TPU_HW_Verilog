module GEMM #(
    // Parameter
    parameter DATA_WIDTH = 8,
    parameter PSUM_WIDTH = 32,
    parameter PE_SIZE = 4,
    
    ) 
    (
    // Port
    input clk,
    input rst_n



    );

endmodule
