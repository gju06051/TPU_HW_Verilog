module PE #(
    // parameter
    parameter DATA_WIDTH = 8,
    parameter IF_ROW_WIDTH = 15,
    parameter FILTER_ROW_WIDTH = 3
    )
    (
    // port
    
    );

    localparam PSUM_WIDTH = IF_ROW_WIDTH - FILTER_ROW_WIDTH - 1;





endmodule