module PE #(
    // parameter
    // FILL HERE //
    )
    (
    // port
    // FILL HERE //
    );




endmodule