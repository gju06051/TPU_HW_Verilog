module Systolic_Array #(
    parameter SA_WIDTH      = 4,
    parameter FIFO_DEPTH    = 4,
    parameter DATA_WIDTH    = 8,
    parameter PSUM_WIDTH    = 32
    )
    (

    );
    
endmodule