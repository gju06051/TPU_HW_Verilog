module eight_bit_multiplier(
    input   [7:0]   A,
    input   [7:0]   B,
    output  [16:0]  Product
);
    wire    [8:0]   pp_1 = {1'b1, !(A[7] && B[0]), (A[6] && B[0]), (A[5] && B[0]), (A[4] && B[0]), (A[3] && B[0]), (A[2] && B[0]), (A[1] && B[0]), (A[0] && B[0])};
    wire    [7:0]   pp_2 = {!(A[7] && B[1]), (A[6] && B[1]), (A[5] && B[1]), (A[4] && B[1]), (A[3] && B[1]), (A[2] && B[1]), (A[1] && B[1]), (A[0] && B[1])};
    wire    [7:0]   pp_3 = {!(A[7] && B[2]), (A[6] && B[2]), (A[5] && B[2]), (A[4] && B[2]), (A[3] && B[2]), (A[2] && B[2]), (A[1] && B[2]), (A[0] && B[2])};
    wire    [7:0]   pp_4 = {!(A[7] && B[3]), (A[6] && B[3]), (A[5] && B[3]), (A[4] && B[3]), (A[3] && B[3]), (A[2] && B[3]), (A[1] && B[3]), (A[0] && B[3])};
    wire    [7:0]   pp_5 = {!(A[7] && B[4]), (A[6] && B[4]), (A[5] && B[4]), (A[4] && B[4]), (A[3] && B[4]), (A[2] && B[4]), (A[1] && B[4]), (A[0] && B[4])};
    wire    [7:0]   pp_6 = {!(A[7] && B[5]), (A[6] && B[5]), (A[5] && B[5]), (A[4] && B[5]), (A[3] && B[5]), (A[2] && B[5]), (A[1] && B[5]), (A[0] && B[5])};
    wire    [7:0]   pp_7 = {!(A[7] && B[6]), (A[6] && B[6]), (A[5] && B[6]), (A[4] && B[6]), (A[3] && B[6]), (A[2] && B[6]), (A[1] && B[6]), (A[0] && B[6])};
    wire    [8:0]   pp_8 = {1'b1, (A[7] && B[7]), !(A[6] && B[7]), !(A[5] && B[7]), !(A[4] && B[7]), !(A[3] && B[7]), !(A[2] && B[7]), !(A[1] && B[7]), !(A[0] && B[7])};

    Exact_4_to_2_Comp EX_1
endmodule